module bcd7seg(
        input  [3:0] b,
        output reg [7:0] h
    );

    //  --0--
    //  |   |
    //  5   1
    //  |-6-|
    //  4   2
    //  |   |
    //  --3--

    always @(b) begin
        case (b)
            4'd0 :
                h = 8'b0000_0011;
            4'd1 :
                h = 8'b1001_1111;
            4'd2 :
                h = 8'b0010_0101;
            4'd3 :
                h = 8'b0000_1101;
            4'd4 :
                h = 8'b1001_1001;
            4'd5 :
                h = 8'b0100_1001;
            4'd6 :
                h = 8'b0100_0001;
            4'd7 :
                h = 8'b0001_1111;
            4'd8 :
                h = 8'b0000_0001;
            4'd9 :
                h = 8'b0000_1001;
            4'd10: // A
                h = 8'b0001_0001;
            4'd11: // b
                h = 8'b0100_0001;
            4'd12: // C
                h = 8'b0110_0011;
            4'd13: // d
                h = 8'b1000_0101;
            4'd14: // E
                h = 8'b0110_0001;
            4'd15: // F
                h = 8'b0111_0001;
            default h = 8'b00000000;
        endcase
    end


endmodule
